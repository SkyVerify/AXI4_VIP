package env_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	import axi_utils_pkg::*;
	import axi_agent_pkg::*;

	`include "axi_env_config.svh"
	`include "axi_scoreboard.svh"
	`include "axi_env.svh"

endpackage : env_pkg
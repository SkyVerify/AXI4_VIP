`timescale 1ns/100ps
`define CYCLE 4 // 250MHz 
`define TDRIVE #(0.2*`CYCLE) // set drive time at 20% of cycle